module FSM
(
    input   wire                DATA_VALID                              ,
    input   wire                PAR_EN                                  ,
    input   wire                ser_done                                ,
    input   wire                CLK                                     ,
    input   wire                RST                                     ,

    output  reg                 ser_en                                  ,
    output  reg     [1:0]       mux_sel                                 ,
    output  reg                 Busy
);

/********************************************************************************************/
/********************************************************************************************/

    reg             [4:0]	    current_state							;
    reg             [4:0]	    next_state								;

/********************************************************************************************/
/********************************************************************************************/

    localparam	s0 = 4'b0001											,
                s1 = 4'b0010											,
                s2 = 4'b0100											,
                s3 = 4'b1000											;

/********************************************************************************************/
/********************************************************************************************/

    always@(posedge CLK or negedge RST)
            begin
            
                if (!RST)
                
                    next_state 		<= 	s0								;
                
                else
                
                    current_state 	<= 	next_state 						;
            
            end

/********************************************************************************************/
/********************************************************************************************/

    always@(*)
        begin

            case(current_state)
            
                s0:
                    begin

                        ser_en  = 1'b0                                  ;              
                        mux_sel = 2'b01                                 ;             
                        Busy    = 1'b0                                  ;

                        if(DATA_VALID)      

                            next_state = s1                             ;

                        else        

                            next_state = s0                             ;    

                    end     

/********************************************************************************************/
/********************************************************************************************/

                s1:     
                    begin       

                        ser_en  = 1'b1                                  ;              
                        mux_sel = 2'b00                                 ;             
                        Busy    = 1'b1                                  ;                    
                        
                        next_state = s2                                 ;
                        

                    end

/********************************************************************************************/
/********************************************************************************************/

                s2:
                    begin

                        ser_en  = 1'b1                                  ;              
                        mux_sel = 2'b10                                 ;             
                        Busy    = 1'b1                                  ;

                        if(ser_done)        
                            begin
                            
                                ser_en  = 1'b0                          ; 

                                if(PAR_EN)

                                    next_state = s3                     ;
                                
                                else        
                                
                                    next_state = s0                     ;
                            end
                        else        

                            next_state = s2                             ;    

                    end  

/********************************************************************************************/
/********************************************************************************************/

                s3:     
                    begin       

                        ser_en  = 1'b0                                  ;              
                        mux_sel = 2'b11                                 ;             
                        Busy    = 1'b1                                  ;

                        next_state = s0                                 ;

                    end  

/********************************************************************************************/
/********************************************************************************************/

                default: next_state = s0						        ;

            endcase

        end

endmodule