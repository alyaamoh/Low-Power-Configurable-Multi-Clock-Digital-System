/********************************************************************************************/
/********************************************************************************************/
/**************************		Author: Alyaa Mohamed    ************************************/
/**************************		Module: ClkDiv	         ************************************/
/********************************************************************************************/
/********************************************************************************************/

module ClkDiv #(parameter WIDTH = 3)
(
    input   wire                    i_ref_clk                                       ,
    input   wire                    i_rst_n                                         ,
    input   wire                    i_clk_en                                        ,
    input   wire  [WIDTH-1:0]       i_div_ratio                                     ,

    output  wire                    o_div_clk
);

/*****************************************************************************************/
/*****************************************************************************************/

    reg           [WIDTH-1:0]       counter                                         ;
    reg                             clk_div                                         ;

/*****************************************************************************************/
/*****************************************************************************************/

    always@(posedge i_ref_clk or negedge i_rst_n)
        begin
            if(!i_rst_n)

                counter   <= 'b0                                                    ;

            else if(i_clk_en)
            
                counter <= (counter == (i_div_ratio-1) ) ? 'b0 : (counter + 'b1)    ;
        
        end

/*****************************************************************************************/
/*****************************************************************************************/

    always @(posedge i_ref_clk or negedge i_rst_n)
        begin

            if(!i_rst_n)
             
                clk_div <= 'b0                                                      ;
            
            else if(i_clk_en)
                    
                clk_div <= (counter < (i_div_ratio/2) ) ?  1'b1 : 1'b0              ; 

        end
   
/*****************************************************************************************/
/*****************************************************************************************/

    assign o_div_clk = (i_clk_en) ? clk_div : i_ref_clk                             ;
    
endmodule