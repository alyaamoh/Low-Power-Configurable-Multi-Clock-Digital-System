/********************************************************************************************/
/********************************************************************************************/
/**************************		Author: Alyaa Mohamed      **********************************/
/**************************		Module: Data_Sync_tb	   **********************************/
/********************************************************************************************/
/********************************************************************************************/
`timescale 1ns/1ps

module Data_Sync_tb()                                                   ;

    parameter 				        NUM_STAGES_tb   = 2 			    ;
    parameter                       BUS_WIDTH_tb    = 8                 ;

/********************************************************************************/
/****************************Internal Signals************************************/

    reg         [BUS_WIDTH_tb-1:0]  Unsync_bus_tb                       ;
    reg                             bus_enable_tb                       ;
    reg                             RST_tb                              ;
    reg                             CLK_tb                              ;

    wire                            enable_pulse_tb                     ;
    wire        [BUS_WIDTH_tb-1:0]  Sync_bus_tb                         ;

/********************************************************************************/
/**************************Clock Period******************************************/

    localparam                      CLK_PERIOD      = 100               ;

/********************************************************************************/
/********************************************************************************/

    initial
        begin
        
            $dumpfile("Data_Sync_tb.vcd") 				                ;
            $dumpvars 									                ;

            Unsync_bus_tb   = 'b0                                       ;
            bus_enable_tb   = 'b0                                       ;
            RST_tb          = 'b0                                       ;
            CLK_tb          = 'b0                                       ;

/********************************************************************************/
/********************************************************************************/

            #(CLK_PERIOD*0.7)
            RST_tb          = 'b1                                       ;
            Unsync_bus_tb   = 8'b11001010                               ;
            bus_enable_tb   = 'b0                                       ;

/********************************************************************************/
/******************************Test Cases****************************************/

            #(CLK_PERIOD*0.3)
            bus_enable_tb   = 'b1                                       ;

            #(CLK_PERIOD*1)
            $display ("\n\nTEST CASE 0")				                ;

            if ((Sync_bus_tb == 'b0) && (enable_pulse_tb == 0))
            
                $display ("\nPassed\n")					                ;

            else
                
                $display ("\nFailed\n")					                ;

/********************************************************************************/
/********************************************************************************/

             #(CLK_PERIOD*2)
            $display ("\n\nTEST CASE 1")				                ;

            if ((Sync_bus_tb == 8'b11001010) && (enable_pulse_tb == 1))
            
                $display ("\nPassed\n")					                ;

            else
                
                $display ("\nFailed\n")					                ;

/********************************************************************************/
/********************************************************************************/

            #(CLK_PERIOD*10)
            $finish										                ;
        end    

/********************************************************************************/
/***************************Clock Generator**************************************/

    always #(CLK_PERIOD*0.5) CLK_tb = !CLK_tb			                ;

/********************************************************************************/
/***********************Instantiation Of The Module******************************/

    Data_Sync #(.NUM_STAGES(NUM_STAGES_tb),.BUS_WIDTH(BUS_WIDTH_tb))
    DUT
    (
        .Unsync_bus(Unsync_bus_tb)                                      ,
        .bus_enable(bus_enable_tb)                                      ,
        .RST(RST_tb)                                                    ,
        .CLK(CLK_tb)                                                    ,

        .enable_pulse(enable_pulse_tb)                                  ,
        .Sync_bus(Sync_bus_tb)                          
    );

endmodule