module FSM
(
    input   wire                DATA_VALID                              ,
    input   wire                PAR_EN                                  ,
    input   wire                ser_done                                ,
    input   wire                CLK                                     ,
    input   wire                RST                                     ,

    output  reg                 ser_en                                  ,
    output  reg     [1:0]       mux_sel                                 ,
    output  reg                 Busy
);

/********************************************************************************************/
/********************************************************************************************/

    reg             [4:0]	    current_state							;
    reg             [4:0]	    next_state								;

/********************************************************************************************/
/********************************************************************************************/

    localparam	IDLE   = 4'b0001									    ,
                Start  = 4'b0010									    ,
                DATA   = 4'b0100									    ,
                Parity = 4'b1000									    ;

/********************************************************************************************/
/********************************************************************************************/

    always@(posedge CLK or negedge RST)
            begin
            
                if (!RST)
                
                    next_state 		<= 	IDLE							;
                
                else
                
                    current_state 	<= 	next_state 						;
            
            end

/********************************************************************************************/
/********************************************************************************************/

    always@(*)
        begin

            case(current_state)
            
                IDLE:
                    begin

                        if(DATA_VALID)      

                            next_state = Start                          ;

                        else        

                            next_state = IDLE                           ;    

                    end     

/********************************************************************************************/
/********************************************************************************************/

                Start:     
                    begin       

                        next_state = DATA                               ;
                        
                    end

/********************************************************************************************/
/********************************************************************************************/

                DATA:
                    begin

                        if(ser_done)        
                            begin

                                if(PAR_EN)

                                    next_state = Parity                 ;
                                
                                else        
                                
                                    next_state = IDLE                   ;

                            end
                        else        

                            next_state = DATA                           ;    

                    end  

/********************************************************************************************/
/********************************************************************************************/

                Parity:     
                    begin       

                        next_state = IDLE                               ;

                    end  

/********************************************************************************************/
/********************************************************************************************/

                default: next_state = IDLE						        ;

            endcase

        end

/********************************************************************************************/
/********************************************************************************************/

    always@(*)
        begin
            ser_en  = 1'b0                                              ;              
            mux_sel = 2'b01                                             ;             
            Busy    = 1'b0                                              ;

            case(current_state)
            
                IDLE:
                    begin

                        ser_en  = 1'b0                                  ;              
                        mux_sel = 2'b01                                 ;             
                        Busy    = 1'b0                                  ;

                    end     

/********************************************************************************************/
/********************************************************************************************/

                Start:     
                    begin       

                        ser_en  = 1'b1                                  ;              
                        mux_sel = 2'b00                                 ;             
                        Busy    = 1'b1                                  ;                                            

                    end

/********************************************************************************************/
/********************************************************************************************/

                DATA:
                    begin

                        ser_en  = 1'b1                                  ;              
                        mux_sel = 2'b10                                 ;             
                        Busy    = 1'b1                                  ;

                        if(ser_done)        
                            
                            ser_en  = 1'b0                              ; 

                    end  

/********************************************************************************************/
/********************************************************************************************/

                Parity:     
                    begin       

                        ser_en  = 1'b0                                  ;              
                        mux_sel = 2'b11                                 ;             
                        Busy    = 1'b1                                  ;

                    end  

/********************************************************************************************/
/********************************************************************************************/

                default:
                    begin

                        ser_en  = 1'b0                                  ;              
                        mux_sel = 2'b01                                 ;             
                        Busy    = 1'b0                                  ;
                    
                    end 

            endcase

        end
endmodule