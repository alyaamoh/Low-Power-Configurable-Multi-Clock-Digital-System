/********************************************************************************************/
/********************************************************************************************/
/**************************		Author: Alyaa Mohamed    ************************************/
/**************************		Module: UART_RX_tb       ************************************/
/********************************************************************************************/
/********************************************************************************************/

`timescale 1ns/1ps

module UART_RX_tb();

    parameter   DATA_WIDTH_tb     = 8                           ,
                PRESCALE_WIDTH_tb = 6                           ;

/********************************************************************************************/
/********************************************************************************************/

    reg                                 PAR_EN_tb               ;
    reg                                 RX_IN_tb                ;
    reg  [PRESCALE_WIDTH_tb - 1 : 0]    Prescale_tb             ;
    reg                                 PAR_TYP_tb              ;
    reg                                 RX_CLK_tb               ;
    reg                                 RST_tb                  ;

    wire   [DATA_WIDTH_tb - 1 : 0]      P_DATA_tb               ;
    wire                                data_valid_tb           ;

/********************************************************************************************/
/********************************************************************************************/

    reg                                 TX_CLK_tb               ;
    reg                                 Data_Stimulus_En        ;
    reg   [PRESCALE_WIDTH_tb-1:0]       count                   ;

    reg   [21:0]                        Data = 22'b10011111010_10010101010 ;

/********************************************************************************************/
/********************************************************************************************/

    localparam              CLK_PERIOD      = 100               ;

/********************************************************************************************/
/********************************************************************************************/

    initial
            begin
                
                $dumpfile("UART_RX_tb.vcd") 		            ;
                $dumpvars 							            ;

                PAR_EN_tb        = 'b0                          ;
                RX_IN_tb         = 'b1                          ;
                Prescale_tb      = 'b0                          ;
                PAR_TYP_tb       = 'b0                          ;
                RX_CLK_tb        = 'b1                          ;
                RST_tb           = 'b0                          ;
                TX_CLK_tb        = 'b0                          ;
                Data_Stimulus_En = 'b0                          ;
                count            = 'b0                          ;           

                #CLK_PERIOD
                PAR_EN_tb        = 'b1                          ;
                Prescale_tb      = 'd8                          ;
                PAR_TYP_tb       = 'b0                          ;
                RST_tb           = 'b1                          ;

                #(CLK_PERIOD*10)
                Data_Stimulus_En = 'b1                          ;

                #(CLK_PERIOD*4000)
                $finish                                         ;

            end

/********************************************************************************************/
/********************************************************************************************/

    always @ (posedge TX_CLK_tb)
        begin

            if(Data_Stimulus_En && count < 'd22 )
                begin

                    RX_IN_tb <= Data[count]                     ;
                    count <= count + 'b1                        ;

                end	
            else

                RX_IN_tb <= 'b1                                 ;  

        end

/********************************************************************************************/
/********************************************************************************************/

    always@(posedge RX_CLK_tb)
        begin

            if(data_valid_tb)

                $display("\n\nThe Data is : %b\n\n",P_DATA_tb)  ;

        end

/********************************************************************************************/
/********************************************************************************************/

    always #CLK_PERIOD      RX_CLK_tb = ~RX_CLK_tb              ;

    always #(CLK_PERIOD*8)  TX_CLK_tb = ~TX_CLK_tb              ;

/********************************************************************************************/
/********************************************************************************************/

    UART_RX #(.DATA_WIDTH(DATA_WIDTH_tb), .PRESCALE_WIDTH(PRESCALE_WIDTH_tb)) 
    DUT
    (
        .PAR_EN(PAR_EN_tb)                                      ,
        .RX_IN(RX_IN_tb)                                        ,
        .Prescale(Prescale_tb)                                  ,
        .PAR_TYP(PAR_TYP_tb)                                    ,
        .CLK(RX_CLK_tb)                                         ,
        .RST(RST_tb)                                            ,

        .P_DATA(P_DATA_tb)                                      ,
        .data_valid(data_valid_tb)
    );

endmodule