/********************************************************************************************/
/********************************************************************************************/
/**************************		Author: Alyaa Mohamed      **********************************/
/**************************		Module: UART_TX_tb	       **********************************/
/********************************************************************************************/
/********************************************************************************************/
`timescale 1ns/1ps

module UART_TX_tb ()                                                    ;
    parameter                   WIDTH = 8                               ;

    reg         [WIDTH-1:0]     P_DATA_tb                               ;
    reg                         DATA_VALID_tb                           ;
    reg                         PAR_EN_tb                               ;
    reg                         PAR_TYP_tb                              ;
    reg                         CLK_tb                                  ;
    reg                         RST_tb                                  ;

    wire                        TX_OUT_tb                               ;
    wire                        Busy_tb                                 ;

/********************************************************************************************/
/********************************************************************************************/

    integer                     i                                       ;
    reg         [10:0]          out                                     ;

/********************************************************************************************/
/********************************************************************************************/

    localparam                  CLK_PERIOD = 5                          ;

/********************************************************************************************/
/********************************************************************************************/

    initial 
        begin

            $dumpfile("UART_TX_tb.vcd")                                 ;
            $dumpvars 										            ;

            P_DATA_tb       = 'b0                                       ;
            DATA_VALID_tb   = 'b0                                       ;
            PAR_EN_tb       = 'b0                                       ;
            PAR_TYP_tb      = 'b0                                       ;
            CLK_tb          = 'b0                                       ;

/********************************************************************************************/
/********************************************************************************************/

            #(CLK_PERIOD*0.3)
            RST_tb 		    = 1		                                    ;	

            #(CLK_PERIOD*0.4)
            RST_tb 		    = 0		                                    ;						

            #(CLK_PERIOD*0.3)
            RST_tb 		    = 1								            ;

            $monitor ("Busy Flag %d", Busy_tb)                          ;

/********************************************************************************************/
/******************************************Test 1********************************************/
/**************************************with even parity**************************************/

            #CLK_PERIOD
            P_DATA_tb       = 8'b11001011                               ;
            DATA_VALID_tb   = 'b1                                       ;
            PAR_EN_tb       = 'b1                                       ;
            PAR_TYP_tb      = 'b0                                       ;

            $display ("\n\nTEST CASE 1")					            ;
            #CLK_PERIOD

            for(i=0;i<12;i=i+1)
                begin

                    #CLK_PERIOD
                    DATA_VALID_tb   = 'b0                               ;
                    out[i]          = TX_OUT_tb                         ;

                end

            #(CLK_PERIOD*4)

            if ( out == 11'b11110010110 )				
                
                $display ("\nPassed\n")							        ;

            else

                $display ("\nFailed\n")							        ;

/********************************************************************************************/
/******************************************Test 2********************************************/
/**************************************with odd parity***************************************/

            #CLK_PERIOD
            P_DATA_tb       = 8'b11001011                               ;
            DATA_VALID_tb   = 'b1                                       ;
            PAR_EN_tb       = 'b1                                       ;
            PAR_TYP_tb      = 'b1                                       ;

            $display ("\n\nTEST CASE 2")					            ;
            #CLK_PERIOD

            for(i=0;i<12;i=i+1)
                begin

                    #CLK_PERIOD
                    DATA_VALID_tb   = 'b0                               ;
                    out[i]          = TX_OUT_tb                         ;

                end

            #(CLK_PERIOD*4)

            if ( out == 11'b10110010110 )				
                
                $display ("\nPassed\n")							        ;

            else

                $display ("\nFailed\n")							        ;

/********************************************************************************************/
/******************************************Test 3********************************************/
/**************************************with no parity****************************************/

            #CLK_PERIOD
            P_DATA_tb       = 8'b11001011                               ;
            DATA_VALID_tb   = 'b1                                       ;
            PAR_EN_tb       = 'b0                                       ;
            PAR_TYP_tb      = 'b0                                       ;

            $display ("\n\nTEST CASE 3")					            ;
            #CLK_PERIOD

            for(i=0;i<12;i=i+1)
                begin

                    #CLK_PERIOD
                    DATA_VALID_tb   = 'b0                               ;
                    out[i]          = TX_OUT_tb                         ;

                end

            #(CLK_PERIOD*4)

            if ( out == 11'b11110010110 )				
                
                $display ("\nPassed\n")							        ;

            else

                $display ("\nFailed\n")							        ;


            #(CLK_PERIOD*10)
            $finish	                                                    ;

        end

/********************************************************************************************/
/********************************************************************************************/

    always #(CLK_PERIOD*0.5) CLK_tb = !CLK_tb					        ;

/********************************************************************************************/
/********************************************************************************************/

    UART_TX #( .WIDTH(WIDTH) )
    DUT
    (
        .P_DATA(P_DATA_tb)                                              ,
        .DATA_VALID(DATA_VALID_tb)                                      ,
        .PAR_EN(PAR_EN_tb)                                              ,
        .PAR_TYP(PAR_TYP_tb)                                            ,
        .CLK(CLK_tb)                                                    ,
        .RST(RST_tb)                                                    ,

        .TX_OUT(TX_OUT_tb)                                              ,
        .Busy(Busy_tb)
    );

endmodule