/********************************************************************************************/
/********************************************************************************************/
/**************************		Author: Alyaa Mohamed    ************************************/
/**************************		Module: ClkDiv_tb	     ************************************/
/********************************************************************************************/
/********************************************************************************************/

`timescale 1ns/1ps

module ClkDiv_tb();

    parameter               WIDTH_tb        = 3                         ;

/*****************************************************************************************/
/********************************Internal Signals*****************************************/

    reg                     i_ref_clk_tb                                ;
    reg                     i_rst_n_tb                                  ;
    reg                     i_clk_en_tb                                 ;
    reg  [WIDTH_tb-1:0]     i_div_ratio_tb                              ;

    wire                     o_div_clk_tb                               ;

/*****************************************************************************************/
/*******************************Clock Period**********************************************/

    localparam              CLK_PERIOD      = 100                       ;

/*****************************************************************************************/
/*****************************************************************************************/

    initial
        begin
            
            $dumpfile("ClkDiv_tb.vcd") 				                    ;
            $dumpvars 									                ;

            i_ref_clk_tb    = 'b0                                       ;
            i_rst_n_tb      = 'b0                                       ;
            i_clk_en_tb     = 'b0                                       ;
            i_div_ratio_tb  = 'b0                                       ;

/*****************************************************************************************/
/********************Check Any Changes Happens to The Both Clocks*************************/

            $monitor("Ref clk=%b,Div clk=%b",i_ref_clk_tb,o_div_clk_tb) ;

/*****************************************************************************************/
/*****************************************************************************************/

            #CLK_PERIOD
            i_rst_n_tb      = 'b1                                       ;
            i_div_ratio_tb  = 'b100                                     ;

            #(CLK_PERIOD*3)
            i_clk_en_tb     = 'b1                                       ;

/*****************************************************************************************/
/******************************Clock Divided By 4*****************************************/

            $display ("\n\nDivision by 4\n\n");
            #(CLK_PERIOD*8)

/*****************************************************************************************/
/*************************Reset to move to the next case**********************************/

            i_rst_n_tb      = 'b0                                       ;
            i_div_ratio_tb  = 'b101                                     ;        

            #CLK_PERIOD
            i_rst_n_tb      = 'b1                                       ;

/*****************************************************************************************/
/*****************************Clock Divided By 4******************************************/

            $display ("\n\nDivision by 5\n\n")                          ;
            #(CLK_PERIOD*8)

            $finish	                                                    ;

            end

/*****************************************************************************************/
/*******************************Clock Generator*******************************************/

    always #(CLK_PERIOD*0.5) i_ref_clk_tb = !i_ref_clk_tb			    ;

/*****************************************************************************************/
/**************************Instantiation Of The Module************************************/

    ClkDiv #(.WIDTH(WIDTH_tb))
    DUT
    (
        .i_ref_clk(i_ref_clk_tb)                                        ,
        .i_rst_n(i_rst_n_tb)                                            ,
        .i_clk_en(i_clk_en_tb)                                          ,
        .i_div_ratio(i_div_ratio_tb)                                    ,

        .o_div_clk(o_div_clk_tb)
    );

endmodule