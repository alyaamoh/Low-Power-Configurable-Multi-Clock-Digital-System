module edge_bit_counter
(
    input   wire            enable                                  ,
    input   wire    [5:0]   Prescale                                ,
    input   wire            CLK                                     ,
    input   wire            RST                                     ,

    output  reg     [4:0]   bit_cnt                                 ,
    output  reg     [5:0]   edge_cnt
);

/********************************************************************************************/
/********************************************************************************************/

    wire                    edge_cnt_done                           ;

/********************************************************************************************/
/********************************************************************************************/

    assign edge_cnt_done = (edge_cnt == Prescale) ? 1'b1 : 1'b0     ; 

/********************************************************************************************/
/********************************************************************************************/

    always@(posedge CLK or negedge RST)
        begin

            if(!RST)

                edge_cnt <= 'b0                                     ;
                
            else if( (enable) && (!edge_cnt_done) )
                
                edge_cnt <= edge_cnt + 'd1                          ;

            else

                edge_cnt <= 'b0                                     ;

        end

/********************************************************************************************/
/********************************************************************************************/

    always@(posedge CLK or negedge RST)
        begin

            if(!RST)

                bit_cnt <= 'b0                                      ;
                
            else if( (enable) && (edge_cnt_done) )
                
                bit_cnt <= bit_cnt + 'd1                            ;

            else

                edge_cnt <= 'b0                                     ;

        end    

endmodule