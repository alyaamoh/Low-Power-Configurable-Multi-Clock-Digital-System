/********************************************************************************************/
/********************************************************************************************/
/**************************		Author: Alyaa Mohamed      **********************************/
/**************************		Module: RST_Sync_tb	       **********************************/
/********************************************************************************************/
/********************************************************************************************/
`timescale 1ns/1ps

module RST_Sync_tb()                                            ;

    parameter 				NUM_STAGES_tb   = 2 			    ;

/********************************************************************************/
/*****************************Internal Signals***********************************/

    reg                     RST_tb                              ;
    reg                     CLK_tb                              ;

    wire                    Sync_RST_tb                         ;

/********************************************************************************/
/******************************Clock Period**************************************/

    localparam              CLK_PERIOD      = 100               ;

/********************************************************************************/
/********************************************************************************/

    initial
        begin
        
            $dumpfile("RST_Sync_tb.vcd") 				        ;
            $dumpvars 									        ;

            CLK_tb = 'b0                                        ;

/********************************************************************************/
/******************************Test Cases****************************************/

            RST_tb = 1'b1                                       ;
            #(CLK_PERIOD*3) 

            $display ("\n\nTEST CASE 0")				        ;

            if (Sync_RST_tb == 1 )
            
                $display ("\nPassed\n")					        ;

            else
                
                $display ("\nFailed\n")					        ;


/********************************************************************************/
/********************************************************************************/

            #(CLK_PERIOD*0.7)
            RST_tb = 1'b0                                       ;

            #(CLK_PERIOD*0.4)
            RST_tb = 1'b1                                       ;

            #(CLK_PERIOD*0.9)
            $display ("\n\nTEST CASE 1")				        ;

            if (Sync_RST_tb == 0 )
            
                $display ("\nPassed\n")					        ;

            else
                
                $display ("\nFailed\n")					        ;

/********************************************************************************/
/********************************************************************************/

            #(CLK_PERIOD*2) 

            $display ("\n\nTEST CASE 2")				        ;

            if (Sync_RST_tb == 1 )
            
                $display ("\nPassed\n")					        ;

            else
                
                $display ("\nFailed\n")					        ;    

            #(CLK_PERIOD*10)
            $finish										        ;
        end

/********************************************************************************/
/****************************Clock Generator*************************************/

    always #(CLK_PERIOD*0.5) CLK_tb = !CLK_tb			        ;

/********************************************************************************/
/**********************Instantiation Of The Module*******************************/

    RST_Sync #(.NUM_STAGES(NUM_STAGES_tb))
    DUT
    (
        .RST(RST_tb)                                            ,
        .CLK(CLK_tb)                                            ,

        .Sync_RST(Sync_RST_tb)    
    );

endmodule
