/********************************************************************************************/
/********************************************************************************************/
/**************************		Author: Alyaa Mohamed    ************************************/
/**************************		Module: BIT_SYNC_tb	     ************************************/
/********************************************************************************************/
/********************************************************************************************/

`timescale 1ns/1ps

module BIT_SYNC_tb()                                                ;

    parameter 				    NUM_STAGES_tb   = 2 			    ;
    parameter                   BUS_WIDTH_tb    = 4                 ;

/********************************************************************************/
/*******************************Internal Signals*********************************/

    reg     [BUS_WIDTH_tb-1:0]  ASYNCH_tb                           ;
    reg                         RST_tb                              ;
    reg                         CLK_tb                              ;

    wire    [BUS_WIDTH_tb-1:0]  SYNC_tb                             ;

/********************************************************************************/
/********************************Clock Period************************************/

    localparam                  CLK_PERIOD      = 100               ;

/********************************************************************************/
/********************************************************************************/

    initial
        begin
        
            $dumpfile("BIT_SYNC_tb.vcd") 				            ;
            $dumpvars 									            ;

            CLK_tb      = 'b0                                       ;
            ASYNCH_tb   = 'b0                                       ;
            RST_tb      = 'b0                                       ;

            #(CLK_PERIOD*0.7)
            RST_tb      = 'b1                                       ;

/********************************************************************************/
/***********************************Test Cases***********************************/

            #(CLK_PERIOD*0.3)
            ASYNCH_tb   = 'b1101                                    ;

            #(CLK_PERIOD*3)
            $display ("\n\nTEST CASE 0")				            ;

            if (SYNC_tb == 'b1101 )
            
                $display ("\nPassed\n")					            ;

            else
                
                $display ("\nFailed\n")					            ;

/********************************************************************************/
/********************************************************************************/

            #(CLK_PERIOD*10)
            $finish										            ;
        end    

/********************************************************************************/
/*****************************Clock Generator************************************/

    always #(CLK_PERIOD*0.5) CLK_tb = !CLK_tb			            ;

/********************************************************************************/
/************************Instantiation Of The Module*****************************/

    BIT_SYNC #(.NUM_STAGES(NUM_STAGES_tb), .BUS_WIDTH(BUS_WIDTH_tb))
    DUT
    (
        .ASYNCH(ASYNCH_tb)                                          ,      								
        .RST(RST_tb)                                                ,   								
        .CLK(CLK_tb)                                                ,   								

        .SYNC(SYNC_tb)
    );

endmodule